module top(a, b, c);
	input [3:0] a, b;
	output [7:0] c;

	assign c = a * b;
endmodule
